
module andgate(
input a,b,
output c
    );
    
 //   assign c = a&b;
    and (c,a,b)
endmodule
