module and_gate(
    input a,
    input b,
    output y
    );
    xor(y,a,b);
endmodule
