module main;
  initial 
      $display("Hello, World");
    end
endmodule
